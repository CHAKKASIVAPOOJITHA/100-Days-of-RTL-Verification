module logic_gates(input a,b,output reg and_gate,or_gate,not_gate,nand_gate,nor_gate,xor_gate,xnor_gate);
  assign and_gate=a&b;
  assign or_gate=a|b;
  assign not_gate=~a;
  assign nand_gate=~(a&b);
  assign nor_gate=~(a|b);
  assign nor_gate=a^b;
  assign xnor_gate=~(a^b);
endmodule
